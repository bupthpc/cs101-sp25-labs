module Synchronizer (
    input  clk,
    input  async_in,
    output sync_out
);

  // TODO: implement this

endmodule
