module SevenSegments (
    input [3:0] in,
    output reg [6:0] out
);
    
    // TODO: implement this

endmodule
