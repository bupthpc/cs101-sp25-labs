module top (
    input CLK100MHZ,
    input BTNU,  // up button for increase counter
    input BTNC,  // center button for reset
    output CA, CB, CC, CD, CE, CF, CG,  // seven segments
    output [7:0] AN
);
  
    // TODO: implement this

endmodule
