// TODO: change these paths if you move the Memory or RegFile instantiation
// to a different module
`define RF_PATH   cpu.rf_inst.mem
`define DMEM_PATH cpu.dmem_inst.mem
`define IMEM_PATH cpu.imem_inst.mem