module EdgeDetector (
    input  clk,
    input  serial_in,
    output edge_detect_pulse
);

  // TODO: implement this

endmodule
