module DisplayController #(
    parameter N = 8
) (
    // TODO: add inputs and outputs
);

  // TODO: implement this

endmodule

