module clk_wiz_0 (
    input clk_in1,
    input reset,
    output clk_out1
);

endmodule