// Don't modify this file
`define RF_PATH   cpu.rf_inst.mem
`define DMEM_PATH cpu.dmem_inst.mem
`define IMEM_PATH cpu.imem_inst.mem