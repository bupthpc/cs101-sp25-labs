module Counter #(
    parameter N = 8  // number of digits
) (
    input clk,
    input rst,
    input en,
    output [N*4-1:0] out
);

  // TODO: implement this

endmodule
